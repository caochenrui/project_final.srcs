module MUSIC(
    input clk,
    input start,
    input rstn,             
    input [2:0]speedup,
    output reg B
);
    reg [24:1]t;
    reg [24:1]total;
    reg clk_out;

    always@(posedge clk,negedge rstn)
        if(~rstn) total<=3125000;
        // else if(speedup==1) total<=3125000;
        else if(speedup==2) total<=1562500;
        else total<=3125000;

    always@(posedge clk,negedge rstn)
        if(~rstn) begin clk_out<=0;t<=total; end
        else if(t==0) begin clk_out<=~clk_out;t<=total; end
        else begin t<=t-1; end


    reg [8:1]state;
    always@(posedge clk_out,negedge rstn)         
        if(~rstn) state<=0;
        else if(start) 
            // if(state!=247)
            state<=state+1;
            // else state<=0;
 
    reg [5:1]m;
    always@(*)
    if(start)
        case(state) 
        0	:m=17;
        1	:m=17;
        2	:m=17;
        3	:m=17;
        4	:m=14;
        5	:m=14;
        6	:m=15;
        7	:m=15;
                 
        8	:m=16;
        9	:m=16;
        10	:m=17;
        11	:m=16;
        12	:m=15;
        13	:m=15;
        14	:m=14;
        15	:m=14;
                 
        16	:m=13;
        17	:m=13;
        18	:m=13;
        19	:m=13;
        20	:m=13;
        21	:m=13;
        22	:m=15;
        23	:m=15;
                 
        24	:m=17;
        25	:m=17;
        26	:m=17;
        27	:m=17;
        28	:m=16;
        29	:m=16;
        30	:m=15;
        31	:m=15;
                 
        32	:m=14;
        33	:m=14;
        34	:m=14;
        35	:m=14;
        36	:m=14;
        37	:m=14;
        38	:m=15;
        39	:m=15;
                 
        40	:m=16;
        41	:m=16;
        42	:m=16;
        43	:m=16;
        44	:m=17;
        45	:m=17;
        46	:m=17;
        47	:m=17;
                 
        48	:m=15;
        49	:m=15;
        50	:m=15;
        51	:m=15;
        52	:m=13;
        53	:m=13;
        54	:m=13;
        55	:m=13;

        56	:m=13;
        57	:m=13;
        58	:m=13;
        59	:m=13;
        60	:m=13;
        61	:m=13;
        62	:m=13;
        63	:m=13;

        64	:m=0;
        65	:m=0;
        66	:m=16;
        67	:m=16;
        68	:m=16;
        69	:m=16;
        70	:m=18;
        71	:m=18;

        72	:m=20;
        73	:m=20;
        74	:m=20;
        75	:m=20;
        76	:m=19;
        77	:m=19;
        78	:m=18;
        79	:m=18;

        80	:m=17;
        81	:m=17;
        82	:m=17;
        83	:m=17;
        84	:m=17;
        85	:m=17;
        86	:m=15;
        87	:m=15;

        88	:m=17;
        89	:m=17;
        90	:m=17;
        91	:m=17;
        92	:m=16;
        93	:m=16;
        94	:m=15;
        95	:m=15;

        96	:m=14;
        97	:m=14;
        98	:m=14;
        99	:m=14;
        100	:m=14;
        101	:m=14;
        102	:m=15;
        103	:m=15;

        104	:m=16;
        105	:m=16;
        106	:m=16;
        107	:m=16;
        108	:m=17;
        109	:m=17;
        110	:m=17;
        111	:m=17;

        112	:m=15;
        113	:m=15;
        114	:m=15;
        115	:m=15;
        116	:m=13;
        117	:m=13;
        118	:m=13;
        119	:m=13;

        120	:m=13;
        121	:m=13;
        122	:m=13;
        123	:m=13;
        124	:m=0;
        125	:m=0;
        126	:m=0;
        127	:m=0;

        128	:m=10;
        129	:m=10;
        130	:m=10;
        131	:m=10;
        132	:m=10;
        133	:m=10;
        134	:m=10;
        135	:m=10;

        136	:m=8;
        137	:m=8;
        138	:m=8;
        139	:m=8;
        140	:m=8;
        141	:m=8;
        142	:m=8;
        143	:m=8;

        144	:m=9;
        145	:m=9;
        146	:m=9;
        147	:m=9;
        148	:m=9;
        149	:m=9;
        150	:m=9;
        151	:m=9;

        152	:m=7;
        153	:m=7;
        154	:m=7;
        155	:m=7;
        156	:m=7;
        157	:m=7;
        158	:m=7;
        159	:m=7;

        160	:m=8;
        161	:m=8;
        162	:m=8;
        163	:m=8;
        164	:m=8;
        165	:m=8;
        166	:m=8;
        167	:m=8;

        168	:m=6;
        169	:m=6;
        170	:m=6;
        171	:m=6;
        172	:m=6;
        173	:m=6;
        174	:m=6;
        175	:m=6;

        176	:m=30;//5.5
        177	:m=30;//5.5
        178	:m=30;//5.5
        179	:m=30;//5.5
        180	:m=30;//5.5
        181	:m=30;//5.5
        182	:m=30;//5.5
        183	:m=30;//5.5

        184	:m=7;
        185	:m=7;
        186	:m=7;
        187	:m=7;
        188	:m=0;
        189	:m=0;
        190	:m=0;
        191	:m=0;

        192	:m=10;
        193	:m=10;
        194	:m=10;
        195	:m=10;
        196	:m=10;
        197	:m=10;
        198	:m=10;
        199	:m=10;

        200	:m=8;
        201	:m=8;
        202	:m=8;
        203	:m=8;
        204	:m=8;
        205	:m=8;
        206	:m=8;
        207	:m=8;

        208	:m=9;
        209	:m=9;
        210	:m=9;
        211	:m=9;
        212	:m=9;
        213	:m=9;
        214	:m=9;
        215	:m=9;

        216	:m=7;
        217	:m=7;
        218	:m=7;
        219	:m=7;
        220	:m=7;
        221	:m=7;
        222	:m=7;
        223	:m=7;
        
        224	:m=8;
        225	:m=8;
        226 :m=8;
        227 :m=8;
        228	:m=10;
        229	:m=10;
        230 :m=10;
        231 :m=10;

        232	:m=13;
        233	:m=13;
        234	:m=13;
        235	:m=13;
        236	:m=13;
        237	:m=13;
        238	:m=13;
        239	:m=13;
        240	:m=31;//12.5
        241	:m=31;//12.5
        242	:m=31;//12.5
        243	:m=31;//12.5
        244	:m=31;//12.5
        245	:m=31;//12.5
        246	:m=31;//12.5
        247	:m=31;//12.5
        248	:m=0;
        249	:m=0;
        250	:m=0;
        251	:m=0;
        252 :m=0;
        253 :m=0;
        254 :m=0;
        255 :m=0;
        default: m=0;
        endcase
    else m=0;

    reg [27:1]q;
    always@(*)
    begin
        case(m)
        0 :q=0;
        1 :q=100000000/261 ; //261.6HZ 低do//10000000
        2 :q=100000000/293 ; //293.7HZ 低ri           
        3 :q=100000000/329 ; //329.6HZ 低mi 
        4 :q=100000000/349 ; //349.2HZ 低fa               
        5 :q=100000000/392 ; //392HZ 低so                  
        6 :q=100000000/440 ; //440HZ 低la              
        7 :q=100000000/499 ; //493.9HZ 低xi  
        8 :q=100000000/523 ; //523.3HZ中do
        9 :q=100000000/587 ; //587.3HZ 中ri          
        10:q=100000000/659 ; //659.3HZ 中mi        
        11:q=100000000/698 ; //698.5HZ 中fa
        12:q=100000000/784 ; //784HZ 中so      
        13:q=100000000/880 ; //880HZ 中la            
        14:q=100000000/998 ; //987.8HZ 中xi
        15:q=100000000/1046; //1045.4HZ 高do      
        16:q=100000000/1174; //1174.7HZ 高ri         
        17:q=100000000/1318; //1318.5HZ 高mi
        18:q=100000000/1396; //1396.3HZ 高fa         
        19:q=100000000/1568; //1568HZ 高so           
        20:q=100000000/1760; //1760HZ 高la              
        21:q=100000000/1976; //1975.5HZ 高xi  
        30:q=100000000/415;  //5.5
        31:q=100000000/831;  //12.5                  
        default:q=0;
        endcase    
    end
 
    reg [27:1]p;
    reg [27:1]tt;
    always@(posedge clk,negedge rstn)      
    begin
        if(~rstn) begin B<=0;p<=0; end
        else begin
            tt<=q;
            if(q==0||tt!=q)
            begin
                if(q==0) begin B<=0; end
                if(tt!=q) begin p<=0; end
            end
            else
            begin 
                if(p==q-1) p<=0;
                else p<=p+1;
                if(p==0) B<=1;
                if(p==q/256) B<=0;//占空比控制音量
            end
        end
    end 

endmodule